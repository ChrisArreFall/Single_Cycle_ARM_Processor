module processorTest();

endmodule