module adderARM#(parameter N = 32)(input logic [N-1:0] A,B,
											 output logic [N-1:0] out);
	assign out = A + B;						 
endmodule 

